`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/07/2025 05:43:27 PM
// Design Name: 
// Module Name: ALU_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ALU_tb();

reg [3:0] sel;
reg [31:0] a, b;
wire [31:0] out;
wire zero;
ALU #(32) alu(.sel(sel), .a(a), .b(b), .out(out), .zero(zero));
initial begin
//Addition (b0010)
sel = 4'b0010;
a = 32'b00000111011001011111011111110011; //124123123 
b = 32'b00000100000000111111001010001111; //67367567 
//result = 191490690
#10 
a = 32'b00000000100110001001011010000000; // 10000000 
b = 32'b11111111011001110110100110000000; // -10000000
//result = 0
#10  //Subtraction
sel = 4'b0110;
a = 32'b00000111011001011111011111110011; //124123123 
b = 32'b00000100000000111111001010001111; //67367567 
//result = 56755556
#10 
a = 32'b00000000100110001001011010000000; // 10000000 
b = 32'b00000000100110001001011010000000; // 10000000 
//result = 0
#10  //Anding
sel = 4'b0000;
a = 32'b00000111011001011111011111110011; //124123123 
b = 32'b00000100000000111111001010001111; //67367567 
//result = 67236483 | 100000000011111001010000011
#10 
a = 32'b11111111111111111111111111111111; //-1 
b = 32'b00000000000000000000000000000000; //0 
//result = 0
#10 
sel = 4'b0001;
a = 32'b00000111011001011111011111110011; //124123123 
b = 32'b00000100000000111111001010001111; //67367567 
//result = 124254207 | 111011001111111011111111111 
#10 
a = 32'b00000000000000000000000000000000; //0 
b = 32'b00000000000000000000000000000000; //0 
//result = 0
#10 
sel = 4'b1111;
//result = 0;

end
endmodule
