`timescale 1ns / 1ps


module InstrMem(
input [5:0] addr, output [31:0] data_out
    );
    reg [31:0] memory[0:63];
    assign data_out = memory[addr];
    initial begin
//        /*
        // testing both stalling and forwatding
        memory[0]=32'b000000000000_00000_010_00001_0000011 ; //lw x1, 0(x0)
        memory[1]=32'b000000000100_00000_010_00010_0000011 ; //lw x2, 4(x0)
        memory[2]=32'b000000001000_00000_010_00011_0000011 ; //lw x3, 8(x0)
        memory[3]=32'b0000000_00010_00001_110_00100_0110011 ; //or x4, x1, x2
        memory[4]=32'b00000000001100100000101001100011; //beq x4, x3, 20
        memory[5]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[6]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[7]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[8]=32'b0000000_00010_00001_000_00011_0110011 ; //add x3, x1, x2
        memory[9]=32'b0000000_00010_00011_000_00101_0110011 ; //add x5, x3, x2
        memory[10]=32'b0000000_00101_00000_010_01100_0100011; //sw x5, 12(x0)
        memory[11]=32'b000000001100_00000_010_00110_0000011 ; //lw x6, 12(x0)
        memory[12]=32'b0000000_00001_00110_111_00111_0110011 ; //and x7, x6, x1
        memory[13]=32'b0100000_00010_00001_000_01000_0110011 ; //sub x8, x1, x2
        memory[14]=32'b0000000_00010_00001_000_00000_0110011 ; //add x0, x1, x2
        memory[15]=32'b0000000_00001_00000_000_01001_0110011 ; //add x9, x0, x1
//        */

/*
        //        Testing for only forwarding hazard
        memory[0]=32'b000000000000_00000_010_00001_0000011 ; //lw x1, 0(x0)
        memory[1]=32'b000000000100_00000_010_00010_0000011 ; //lw x2, 4(x0)
        memory[2]=32'b000000001000_00000_010_00011_0000011 ; //lw x3, 8(x0)
        memory[3]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[4]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[5]=32'b0000000_00010_00001_110_00100_0110011 ; //or x4, x1, x2
        memory[6]=32'b00000000001100100000101001100011; //beq x4, x3, 20
        memory[7]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[8]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[9]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[10]=32'b0000000_00010_00001_000_00011_0110011 ; //add x3, x1, x2
        memory[11]=32'b0000000_00010_00011_000_00101_0110011 ; //add x5, x3, x2
        memory[12]=32'b0000000_00101_00000_010_01100_0100011; //sw x5, 12(x0)
        memory[13]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[14]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[15]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[16]=32'b000000001100_00000_010_00110_0000011 ; //lw x6, 12(x0)
        memory[17]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[18]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[19]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[20]=32'b0000000_00001_00110_111_00111_0110011 ; //and x7, x6, x1
        memory[21]=32'b0100000_00010_00001_000_01000_0110011 ; //sub x8, x1, x2
        memory[22]=32'b0000000_00010_00001_000_00000_0110011 ; //add x0, x1, x2
        memory[23]=32'b0000000_00001_00000_000_01001_0110011 ; //add x9, x0, x1
*/
        /*
        // Remove all possible NOPs without any hazards units to counter
        memory[0]=32'b000000000000_00000_010_00001_0000011 ; //lw x1, 0(x0)
        memory[1]=32'b000000000100_00000_010_00010_0000011 ; //lw x2, 4(x0)
        memory[2]=32'b000000001000_00000_010_00011_0000011 ; //lw x3, 8(x0)
        memory[3]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[4]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[5]=32'b0000000_00010_00001_110_00100_0110011 ; //or x4, x1, x2
        memory[6]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[7]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[8]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[9]=32'b00000010001100100000000001100011; //beq x4, x3, 32
        memory[10]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[11]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[12]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[13]=32'b0000000_00010_00001_000_00011_0110011 ; //add x3, x1, x2
        memory[14]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[15]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[16]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[17]=32'b0000000_00010_00011_000_00101_0110011 ; //add x5, x3, x2
        memory[18]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[19]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[20]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[21]=32'b0000000_00101_00000_010_01100_0100011; //sw x5, 12(x0)
        memory[22]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[23]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[24]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[25]=32'b000000001100_00000_010_00110_0000011 ; //lw x6, 12(x0)
        memory[26]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[27]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[28]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
        memory[29]=32'b0000000_00001_00110_111_00111_0110011 ; //and x7, x6, x1
        memory[30]=32'b0100000_00010_00001_000_01000_0110011 ; //sub x8, x1, x2
        memory[31]=32'b0000000_00010_00001_000_00000_0110011 ; //add x0, x1, x2
        memory[32]=32'b0000000_00001_00000_000_01001_0110011 ; //add x9, x0, x1
        */
        
        
        //No NOPs
        /*
        memory[0]=32'b000000000000_00000_010_00001_0000011 ; //lw x1, 0(x0)
        memory[1]=32'b000000000100_00000_010_00010_0000011 ; //lw x2, 4(x0)
        memory[2]=32'b000000001000_00000_010_00011_0000011 ; //lw x3, 8(x0)
        memory[3]=32'b0000000_00010_00001_110_00100_0110011 ; //or x4, x1, x2
        memory[4]=32'b00000000001100100000010001100011; //beq x4, x3, 8
        memory[5]=32'b0000000_00010_00001_000_00011_0110011 ; //add x3, x1, x2
        memory[6]=32'b0000000_00010_00011_000_00101_0110011 ; //add x5, x3, x2
        memory[7]=32'b0000000_00101_00000_010_01100_0100011; //sw x5, 12(x0)
        memory[8]=32'b000000001100_00000_010_00110_0000011 ; //lw x6, 12(x0)
        memory[9]=32'b0000000_00001_00110_111_00111_0110011 ; //and x7, x6, x1
        memory[10]=32'b0100000_00010_00001_000_01000_0110011 ; //sub x8, x1, x2
        memory[11]=32'b0000000_00010_00001_000_00000_0110011 ; //add x0, x1, x2
        memory[12]=32'b0000000_00001_00000_000_01001_0110011 ; //add x9, x0, x1
        */
        
        //The looping code way back then
        /*
        memory[0]=32'b00000000000000000010000100000011 ; //lw x2, 0(x0)
        memory[1]=32'b00000000010000000010000110000011 ; //lw x3, 4(x0)
        memory[2]=32'b00000000000000000000000010110011 ; //add x1, x0, x0
        memory[3]=32'b00000000001000001000000010110011 ; //add x1, x1, x2
        memory[4]=32'b00000000001100001110001000110011 ; //or x4, x1, x3
        memory[5]=32'b11111110001100100000110011100011 ; //beq x4, x3, -8
        memory[6]=32'b00000000010000000010010000100011 ; //sw x4, 8(x0)
        memory[7]=32'b01000000001100100000001010110011 ; //sub x5, x4, x3
        memory[8]=32'b00000000001000101111001100110011 ; //and x6, x5, x2
        */
    end
    
endmodule
