`timescale 1ns / 1ps

module ImmGen_tb();
reg [31:0] in;
wire [31:0] imm;

ImmGen immediateGenerator(.instr(in), .imm(imm));
initial begin
//For SW and LW
//010011010010 -- 1234
//001100010011 -- 787
//111001011001 -- -423
//110000011000 -- -1000


//Start of LW
in = 32'b01001101001000000000000000010011; // Imm = 1234
#10 
in = 32'b00110001001100000000000000010011; // Imm = 787
#10 
in = 32'b11100101100100000000000000010011; // Imm = -423
#10 
in = 32'b11000001100000000000000000010011; // Imm = -1000 
//Start of SW
#10 
in = 32'b01001100000000000000100100100011; // 1234
#10
in = 32'b00110000000000000000100110100011; // 787
#10 
in = 32'b11100100000000000000110010100011; // -423
#10 
in = 32'b11000000000000000000110000100011; // -1000
//For BEQ
// 1010010001110 = -2930
// 0011110001010 = 1930
//Start of BEQ 
in = 32'b11001000000000000000011101100011; // -2930
#10 
in = 32'b01111000000000000000010101100011; // 1930


end

endmodule
